`include "uvm_pkg.sv"	//for compilation
`include "uvm_macros.svh"
import uvm_pkg::*;		//for making them available
`include "./common/axi_config.sv"
`include "./common/axi_interface.sv"
`include "./top/axi_assertions.sv"
`include "./slave/memory.v"
`include "./common/axi_tx.sv"
`include "./master/axi_seq_lib.sv"
`include "./master/axi_sqr.sv"
`include "./master/axi_driver.sv"
`include "./common/axi_mon.sv"
`include "./master/axi_cov.sv"
`include "./slave/axi_responder.sv"
`include "./master/axi_magent.sv"
`include "./slave/axi_sagent.sv"
`include "./common/axi_sbd_tx_compare.sv"
//`include "./common/axi_sbd_byte_compare.sv"
//`include "./common/axi_sbd_byte_compare_aa.sv"
`include "./top/axi_env.sv"
`include "./top/axi_test.sv"
`include "./top/top.sv"
